module lexer
